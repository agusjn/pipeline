module sra (
    a,
    b,
    o_sra
);
  parameter N = 32;
  input logic [N-1:0] a;
  input logic [N-1:0] b;
  output logic [N-1:0] o_sra;
  logic [N-1:0] o_sra_temp;
  srl srl1 (
      .a(a),
      .b(b),
      .o_srl(o_sra_temp)
  );
  always_comb begin

    if (a[N-1] == 1) begin
      case (b[4:0])
        5'b00000: o_sra <= a;
        5'b00001: o_sra <= {1'b1, a[N-1:1]};
        5'b00010: o_sra <= {2'b11, a[N-1:2]};
        5'b00011: o_sra <= {3'b111, a[N-1:3]};
        5'b00100: o_sra <= {4'b1111, a[N-1:4]};
        5'b00101: o_sra <= {5'b11111, a[N-1:5]};
        5'b00110: o_sra <= {6'b111111, a[N-1:6]};
        5'b00111: o_sra <= {7'b1111111, a[N-1:7]};
        5'b01000: o_sra <= {8'b11111111, a[N-1:8]};
        5'b01001: o_sra <= {9'b111111111, a[N-1:9]};
        5'b01010: o_sra <= {10'b1111111111, a[N-1:10]};
        5'b01011: o_sra <= {11'b11111111111, a[N-1:11]};
        5'b01100: o_sra <= {12'b111111111111, a[N-1:12]};
        5'b01101: o_sra <= {13'b1111111111111, a[N-1:13]};
        5'b01110: o_sra <= {14'b11111111111111, a[N-1:14]};
        5'b01111: o_sra <= {15'b111111111111111, a[N-1:15]};
        5'b10000: o_sra <= {16'b1111111111111111, a[N-1:16]};
        5'b10001: o_sra <= {17'b11111111111111111, a[N-1:17]};
        5'b10010: o_sra <= {18'b111111111111111111, a[N-1:18]};
        5'b10011: o_sra <= {19'b1111111111111111111, a[N-1:19]};
        5'b10100: o_sra <= {20'b11111111111111111111, a[N-1:20]};
        5'b10101: o_sra <= {21'b111111111111111111111, a[N-1:21]};
        5'b10110: o_sra <= {22'b1111111111111111111111, a[N-1:22]};
        5'b10111: o_sra <= {23'b11111111111111111111111, a[N-1:23]};
        5'b11000: o_sra <= {24'b111111111111111111111111, a[N-1:24]};
        5'b11001: o_sra <= {25'b1111111111111111111111111, a[N-1:25]};
        5'b11010: o_sra <= {26'b11111111111111111111111111, a[N-1:26]};
        5'b11011: o_sra <= {27'b111111111111111111111111111, a[N-1:27]};
        5'b11100: o_sra <= {28'b1111111111111111111111111111, a[N-1:28]};
        5'b11101: o_sra <= {29'b11111111111111111111111111111, a[N-1:29]};
        5'b11110: o_sra <= {30'b111111111111111111111111111111, a[N-1:30]};
        5'b11111: o_sra <= {31'b1111111111111111111111111111111, a[N-1:31]};
        default:  o_sra <= 32'h0;
      endcase
    end else begin
      o_sra <= o_sra_temp;
    end
  end
endmodule
